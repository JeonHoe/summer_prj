module testbench();
    
    reg a, b;
    wire sum, c_out;

    halfadd ha1(sum, c_out, a, b);

    initial
    begin
        a = 1'b0; b = 1'b0;
        #10 a = 1'b0; b = 1'b0;
        #10 a = 1'b0; b = 1'b1;
        #10 a = 1'b0; b = 1'b1;
        #10 a = 1'b1; b = 1'b0;
        #10 a = 1'b1; b = 1'b0;
        #10 a = 1'b1; b = 1'b1;
        #10 a = 1'b1; b = 1'b1;
        #10 $stop;
    end

endmodule