module testbench();
    
    reg a, b;
    wire diff, borrow;

    halfsubtract hs1(diff, borrow, a, b);

    initial
    begin
        a = 1'b0; b = 1'b0;
        #10 a = 1'b0; b = 1'b0;
        #10 a = 1'b0; b = 1'b1;
        #10 a = 1'b0; b = 1'b1;
        #10 a = 1'b1; b = 1'b0;
        #10 a = 1'b1; b = 1'b0;
        #10 a = 1'b1; b = 1'b1;
        #10 a = 1'b1; b = 1'b1;
        #10 $stop;
    end

endmodule