`timescale 1ns/1ps
module testbench();
    
    reg a, b;
    wire diff, c_out;

    twos_complement_subtract tcs1 (diff, c_out, a, b);

    initial
    begin
        a = 1'b0; b = 1'b0;
        #10 a=1'b0; b = 1'b1;
        #10 a=1'b1; b = 1'b0;
        #10 a=1'b1; b = 1'b1;
        #10 $stop;

    end

endmodule