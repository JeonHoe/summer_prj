module not_gate(a, out);

    input in;
    output out;

    assign out = ~a;
    
endmodule