module test(input);

    input input0;

endmodule